module map_rom ( input [16:0]	addr,
				 output [11:0]	data
			);

    parameter ADDR_WIDTH = 17;
    parameter DATA_WIDTH =  12;
	logic [ADDR_WIDTH-1:0] addr_reg;
				
	// ROM definition				
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h9DB,
        12'h9DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h9DB,
        12'h9DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h9DB,
        12'h9DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h9DB,
        12'h9DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hEFF,
        12'hEFF,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'hBED,
        12'hBED,
        12'hBED,
        12'hBED,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h8DB,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h9EC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h351,
        12'h351,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h766,
        12'h766,
        12'h766,
        12'h766,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h433,
        12'h433,
        12'h433,
        12'h433,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hAEC,
        12'hAEC,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'hAEC,
        12'hAEC,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h1A6,
        12'h1A6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'hEA7,
        12'h4B8,
        12'h4B8,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'h3A8,
        12'h3A8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'hDEF,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'hDEF,
        12'hDEF,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'hDEB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h8DB,
        12'h8DB,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h4B8,
        12'h4B8,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h4B8,
        12'h4B8,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'h393,
        12'h393,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'hBF8,
        12'hBF8,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h1A6,
        12'h1A6,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h7CA,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h393,
        12'h351,
        12'h351,
        12'h351,
        12'h351,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393,
        12'h8D6,
        12'h8D6,
        12'h393,
        12'h393
    };

	assign data = ROM[addr];

endmodule